module probador (//Entradas
				   output reg clk,      
                   output reg reset_L, 
                   output reg init,    
			       output reg [5:0]  data_in_principal,  
			       output reg push,                    
			       output reg pop_D0,  
			       output reg pop_D1,  

			// output reg [1:0] umbral_MF, 	
	     		// output reg [3:0] umbral_VC0,	
                   	// output reg [3:0] umbral_VC1, 	
	               	// output reg [1:0] umbral_D0, 	
                   	// output reg [1:0] umbral_D1,
                
				   //salidas
				   input [5:0] data_out0, 
			       input [5:0] data_out1, 
			       input active_out,  
				   input idle_out,    
				   input error_out,   
				   input Pausa_MF);
   
// Probador
 initial #0 clk <= 1; // inicia el reloj en 0.
    always
    #1 clk <= ~clk; // el reloj cambia cada ciclo

initial begin
  $dumpfile("test.vcd");
  $dumpvars;

   init <=0 ;
   pop_D0<=0;
   pop_D1<=0;
   push<=0;
   data_in_principal<=0;
   reset_L<=0;

    #2;
	reset_L<=1;

	#1;
    init<=1;
    
    #2;
    init<=0;

    	/////////////////////////////////////////////////
     	//4 PUSH a D0 
     	//2 POP A D0 
     	//2 POP A D1
    	/////////////////////////////////////////////////
	#7; /// 1
    push<=1;
	data_in_principal<=6'b011011; // 0 1 B (VC0,D0,DATA)

	#2;  	/// 2
		data_in_principal<=6'b101101; // 1 0 D
      
   #2;	/// 3;
      		data_in_principal<=6'b000011; // 0 0 3

   #2;		/// 4
      		data_in_principal<=6'b011010; // 0 1 A

	/////////////////////////////////////////////////D
      
   //#2; 
    //  		data_in_principal<=6'b000000; // 0
    
    #2;
		push<=0;	
	//	pop_D0<=1;

	
	//	pop_D0<=1;

	/////////////////////////////////////////////////
/*
	@(posedge clk);		/// 5
		push<=0;
		pop_D0<=0; 
		pop_D1<=1;

	/////////////////////////////////////////////////
     	//2 PUSH a D1
     	//2 PUSH a D0
	//2 PUSH a D0  
    	/////////////////////////////////////////////////
     	@(posedge clk);		/// 6
		push<=1;
		pop_D0<=0; 
		pop_D1<=1;
      		data_in_principal<=6'b111011; // 1 1 B

      	@(posedge clk)		/// 7
		//push<=1;
		pop_D1<=0; 
		data_in_principal<=6'b101011; // 1 1 B

     	@(posedge clk);		/// 8
      		//push<=1;
		pop_D1<=0; 
      		data_in_principal<=6'b001001;// 0 0 9

      	@(posedge clk);		/// 9
      		//push<=1;
      		data_in_principal<=6'b001010;// 0 0 10
	/////////////////////////////////////////////////

	@(posedge clk);		/// 5
		push<=0;    */

#60
   $finish;
end  

   

endmodule 
