
module dual_port_memory # ( parameter DATA_WIDTH= 6, parameter ADDR_WIDTH=8, parameter MEM_SIZE=7 )
(
	input wire						Clock,
	input wire						iWriteEnable,
	input wire [ADDR_WIDTH-1:0]	iReadAddress0,
	input wire [ADDR_WIDTH-1:0]	iWriteAddress,
	input wire [DATA_WIDTH-1:0]		 	iDataIn,
	output reg [DATA_WIDTH-1:0] 		oDataOut0);

reg [DATA_WIDTH-1:0] Ram [MEM_SIZE:0];		

always @(posedge Clock) 
begin 
	
		if (iWriteEnable) 
			Ram[iWriteAddress] <= iDataIn; 
			oDataOut0 <= Ram[iReadAddress0];
		
end 
endmodule

